
module fir (
    input wire clk,
    input wire rst,
    input wire in_valid,
    input logic signed [11:0] in_data,
    output wire in_ready,
    output reg out_valid,
    output logic signed [11:0] out_data,
    input wire out_ready
  );

  real regs [63:0];
  real coefs [0:63] = {
    -6.518263187043542e-19, -7.986557578197472e-04, -0.002095202987291, -0.003667107969085,
    -0.005116643415385, -0.005928729916395, -0.005574799504880, -0.003647417401953,
    4.178988515525191e-18, 0.005140327380087, 0.011118819256345, 0.016883231769783,
    0.021109413050609, 0.022415483902514, 0.019637994970885, 0.012126229259175,
    -8.833912267524514e-18, -0.015685124676703, -0.032911842822594, -0.048841462160068,
    -0.060120550944356, -0.063323725395885, -0.055474603586424, -0.034566931655455,
    1.284346534816169e-17, 0.047150897274960, 0.104087211505337, 0.166488826877401,
    0.228951469309608, 0.285607773393619, 0.330847986488195, 0.360037028336954,
    0.370121787174637, 0.360037028336954, 0.330847986488195, 0.285607773393619,
    0.228951469309608, 0.166488826877401, 0.104087211505337, 0.047150897274960,
    1.284346534816169e-17, -0.034566931655455, -0.055474603586424, -0.063323725395885,
    -0.060120550944356, -0.048841462160068, -0.032911842822594, -0.015685124676703,
    -8.833912267524514e-18, 0.012126229259175, 0.019637994970885, 0.022415483902514, 
    0.021109413050609, 0.016883231769783, 0.011118819256345, 0.005140327380087,
    4.178988515525191e-18, -0.003647417401953, -0.005574799504880, -0.005928729916395,
    -0.005116643415385, -0.003667107969085, -0.002095202987291, -7.986557578197472e-04
  };

  assign out_valid = 1'b1;
  assign in_ready = 1'b1;

  always @(posedge clk) begin
    if(rst) begin
      for(int i =0;i<64;i=i+1) begin
        regs[i] <= 0;
      end
    end
    else begin
      for(int i =0;i<64;i=i+1) begin
        regs[i] <= (i>0) ? (coefs[i]*in_data + regs[i-1]) : coefs[i]*in_data;
      end
      out_data <= regs[63]/4;
    end
  end

endmodule
